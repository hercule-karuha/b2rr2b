WORD_WIDTH 8 BYTE_WIDTH;
typedef 32 WORD_WIDTH;

import "BDPI" function Bit#(n) get(Bit#(WORD_WIDTH) id, Bit#(WORD_WIDTH) cycles, Bit#(WORD_WIDTH) size);
import "BDPI" function Action put(Bit#(WORD_WIDTH) id, Bit#(WORD_WIDTH) cycles, Bit#(n) data, Bit#(WORD_WIDTH) size);


interface RProbe#(type get_t, type put_t);
    method get_t get_data();
    method Action put_data(put_t data);
endinterface

module mkRProbe#(Bit#(WORD_WIDTH) id)(RProbe#(get_t, put_t)) provisos(Bits#(get_t, wid_get), Bits#(put_t, wid_put));
    Bit#(WORD_WIDTH) get_size = fromInteger(valueOf(TDiv#(wid_get, BYTE_WIDTH)));
    Bit#(WORD_WIDTH) put_size = fromInteger(valueOf(TDiv#(wid_put, BYTE_WIDTH)));

    Reg#(Bit#(WORD_WIDTH)) cycles <- mkReg(0);

    rule count;
        cycles <= cycles + 1;
    endrule

    method get_t get_data();
        Bit#(n) data = get(id, cycles, get_size);
        return unpack(data);
    endmethod

    method Action put_data(put_t data);
        let bvec = pack(data);
        put(id, cycles, bvec, put_size);
    endmethod
endmodule