import

module